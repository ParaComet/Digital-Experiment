library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Clk_Generater is
    generic (
        INPUT_CLK : integer := 50_000_000  -- ��ʱ�ӣ�Hz��
    );
    port (
        clk       : in  std_logic;  -- ��ʱ��
        rst       : in  std_logic;  -- �첽��λ������Ч
        clk_1khz  : out std_logic;  -- 1 kHz ʱ�����
        clk_100hz : out std_logic;  -- 100 Hz ʱ�����
        clk_1mhz  : out std_logic   -- 1 MHz ʱ�����
    );
end entity Clk_Generater;

architecture rtl of Clk_Generater is
    -- �����ڼ������� INPUT_CLK ����Ŀ��Ƶ�ʵķ���
    constant HALF_TICKS_1K  : integer := INPUT_CLK / (2 * 1000);
    constant HALF_TICKS_100 : integer := INPUT_CLK / (2 * 100);
    constant HALF_TICKS_1M : integer := INPUT_CLK / (2 * 1_000_000);

    signal cnt1k  : integer := 0;
    signal cnt100 : integer := 0;
    signal cnt1m  : integer := 0;
    signal clk1k_r  : std_logic := '0';
    signal clk100_r : std_logic := '0';
begin

    clk_1khz  <= clk1k_r;
    clk_100hz <= clk100_r;

    process(clk, rst)
    begin
        if rst = '1' then
            cnt1k     <= 0;
            cnt100    <= 0;
            clk1k_r   <= '0';
            clk100_r  <= '0';
        elsif rising_edge(clk) then
            -- 1 MHz ��Ƶ���л�����������
            if cnt1m >= HALF_TICKS_1M - 1 then
                cnt1m <= 0;
            else
                cnt1m <= cnt1m + 1;
            end if;

            -- 1 kHz ��Ƶ���л�����������
            if cnt1k >= HALF_TICKS_1K - 1 then
                cnt1k <= 0;
                clk1k_r <= not clk1k_r;
            else
                cnt1k <= cnt1k + 1;
            end if;

            -- 100 Hz ��Ƶ
            if cnt100 >= HALF_TICKS_100 - 1 then
                cnt100 <= 0;
                clk100_r <= not clk100_r;
            else
                cnt100 <= cnt100 + 1;
            end if;
        end if;
    end process;

end architecture rtl;